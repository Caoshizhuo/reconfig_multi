library verilog;
use verilog.vl_types.all;
entity reconfig_multi_tb is
end reconfig_multi_tb;
